`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2020/02/09 11:45:27
// Design Name:
// Module Name: Tc_PL
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module Tc_PL
#(
parameter TOP0_0	= 3    ,
          TOP0_1	= 7    ,
          TOP0_2	= 2    ,
          TOP0_3	= 12   ,
          TOP0_4	= 4    ,
          ADC0_0  = 14   ,
          ADC0_1  = 56   ,
          LDD0_0  = 32   ,
          CAP0_0  = 4    ,
          CAP0_1  = 2    ,
          AGP0_0	= 3    ,
          AGP0_1	= 2    ,
          AGP0_2	= 1    ,
          AGP0_3	= 3    ,
	        AGP0_4	= 3    ,
	        AGP0_5	= 32   ,
	        AGP0_6	= 8    ,
	        AGP0_7	= 3    ,
	        AGP0_8	= 14   ,
	        AGP0_9	= 32   ,
	        AGP0_10	= 32   ,
	        AGP0_11	= 32   ,
	        AGP0_12	= 18   ,
	        AGP0_13	= 32   ,
	        AGP0_14	= 32   ,
	        AGP0_15	= 6    ,
	        AGP0_16	= 4    ,
	        AGP0_17	= 4    ,
	        AGP0_18	= 5    ,
	        AGP0_19	= 3    ,
	        AGP0_20	= 32   ,
	        AGP0_21	= 6    ,
	        AGP0_22	= 2    ,
	        AGP0_23	= 9    ,
	        AGP0_24	= 8    ,
	        AGP0_25	= 8    ,
	        AGP0_26	= 8    ,
	        AGP0_27	= 16   ,
	        AGP0_28	= 15   ,
	        AGP0_29	= 4    ,
	        AGP0_30	= 2    ,
	        AGP0_31	= 1    ,
	        AGP0_32	= 2    ,
	        AGP0_33	= 1    ,
	        AGP0_34	= 2    ,
	        AGP0_35	= 16
)(
input                     clk125             ,
input                     rst                ,
input                     Gc_adc_of          ,
input      [ADC0_0-1:0]   Gc_adc_data        ,
input                     Gc_cap_mode        ,
output     [TOP0_0-1:0]   Gc_cap_wdis        ,
output     [LDD0_0-1:0]   Gc_cap_plus        ,
output     [TOP0_0-1:0]   Gc_com_wdis        ,
output     [LDD0_0-1:0]   Gc_com_plus        ,
output                    Gc_com_open        ,
output                    Gc_com_close       ,
input      [ADC0_1-1:0]   Gc_merge_data      ,
input                     Gc_mereg_datv      ,
output                    Gc_mereg_datr      ,
output                    Gc_cap_trig        ,
input                     Gc_capr_rdy        ,
input      [TOP0_0-1:0]   Gc_wdis            ,
output     [AGP0_1 -1:0]  gp0_c0	           ,
input                     gp0_c1	           ,
input      [AGP0_2 -1:0]  gp0_c2	           ,
input      [AGP0_3 -1:0]  gp0_c3	           ,
input      [AGP0_4 -1:0]  gp0_c4	           ,
input      [AGP0_5 -1:0]  gp0_c5	           ,
input      [AGP0_6 -1:0]  gp0_c6	           ,
input      [AGP0_7 -1:0]  gp0_c7	           ,
input      [AGP0_8 -1:0]  gp0_c8	           ,
input      [AGP0_9 -1:0]  gp0_c9	           ,
output     [AGP0_10-1:0]  gp0_c10	           ,
output     [AGP0_11-1:0]  gp0_c11	           ,
input      [AGP0_12-1:0]  gp0_c12	           ,
input      [AGP0_12-1:0]  gp0_c13	           ,
input      [AGP0_12-1:0]  gp0_c14	           ,
input      [AGP0_12-1:0]  gp0_c15	           ,
input      [AGP0_13-1:0]  gp0_c16	           ,
input      [AGP0_13-1:0]  gp0_c17	           ,
input      [AGP0_13-1:0]  gp0_c18	           ,
input      [AGP0_13-1:0]  gp0_c19	           ,
input      [AGP0_14-1:0]  gp0_c20	           ,
input      [AGP0_14-1:0]  gp0_c21	           ,
input      [AGP0_14-1:0]  gp0_c22	           ,
input      [AGP0_14-1:0]  gp0_c23	           ,
input      [AGP0_14-1:0]  gp0_c24	           ,
input      [AGP0_14-1:0]  gp0_c25	           ,
input      [AGP0_14-1:0]  gp0_c26	           ,
input      [AGP0_14-1:0]  gp0_c27	           ,
input      [AGP0_15-1:0]  gp0_c28	           ,
input      [AGP0_15-1:0]  gp0_c29	           ,
input      [AGP0_15-1:0]  gp0_c30	           ,
input      [AGP0_15-1:0]  gp0_c31	           ,
input      [AGP0_16-1:0]  gp0_c32	           ,
input      [AGP0_16-1:0]  gp0_c33	           ,
input      [AGP0_16-1:0]  gp0_c34	           ,
input      [AGP0_16-1:0]  gp0_c35	           ,
input      [AGP0_17-1:0]  gp0_d0	           ,
output     [AGP0_18-1:0]  gp0_d1	           ,
input      [AGP0_19-1:0]  gp0_d2	           ,
input      [AGP0_20-1:0]  gp0_d3	           ,
input                     gp0_d4	           ,
input                     gp0_d5	           ,
output     [AGP0_21-1:0]  gp0_b0	           ,
input      [AGP0_22-1:0]  gp0_b1	           ,
input      [AGP0_23-1:0]  gp0_b2	           ,
output     [AGP0_24-1:0]  gp0_b3	           ,
output     [AGP0_25-1:0]  gp0_b4	           ,
output     [AGP0_26-1:0]  gp0_b5	           ,
input      [AGP0_27-1:0]  gp0_b6	           ,
output     [AGP0_28-1:0]  gp0_r0	           ,
input      [AGP0_29-1:0]  gp0_r1	           ,
input      [AGP0_30-1:0]  gp0_r2	           ,
input      [AGP0_31-1:0]  gp0_r3	           ,
output     [AGP0_32-1:0]  gp0_r4	           ,
input      [AGP0_33-1:0]  gp0_r5	           ,
output     [AGP0_34-1:0]  gp0_r6	           ,
input      [AGP0_35-1:0]  gp0_r7             ,
input                     gp0_c0w            ,
input                     gp0_b0w            ,
input                     gp0_b2w  	         ,
input                     gp0_b4r  	         ,
input                     gp0_r7w  	         ,
output                    acp0_tx_en         ,
input                     acp0_tx_rdy        ,
output     [31:0]         acp0_tx_awaddr     ,
output     [2:0]          acp0_tx_awid       ,
output     [63:0]         acp0_tx_wdata      ,
input                     acp0_tx_wdreq      ,
output     [15:0]         IRQ_F2P_0          ,
output                    ADC0_CSN           ,
output                    ADC0_SCK           ,
output                    ADC0_SDI           ,
input                     ADC0_SDO           ,
output                    FDA0_SCK           ,
output                    FDA0_CSN           ,
output                    FDA0_SDI           ,
input                     FDA0_SDO           ,
output                    LDD0_OUTEA         ,
output                    LDD0_DISEA         ,
output                    LDD0_OSCEA         ,
output                    LDD0_OLD2N         ,
output                    LDD0_RDISN         ,
output                    DAC0_SDI           ,
output                    DAC0_SCK           ,
output                    DAC0_CSN           ,
output                    DAC1_SDI           ,
output                    DAC1_SCK           ,
output                    DAC1_CSN           ,
output                    OPA0_10X1          ,
output                    OPA0_10X2          ,
output                    OPA0_OPX1          ,
output                    OPA0_OPX2          ,
output                    APD0_EN            ,
output                    LPL0_CSN           ,
input                     LPL0_SDO           ,
output                    LPL0_SCK           ,
output                    LPL0_SDI           ,
input                     LPL0_LOCK          ,
input                     LPL0_ERR           ,
output                    LPL0_SYNC          ,
input                     TEC0_GOOD          ,
input                     TEC1_GOOD          ,
output     [TOP0_2-1:0]   LED0_L             ,
output     [TOP0_4-1:0]   OPM0_IO
    );

wire        cap_FDA0_SCK   ;
wire        cap_FDA0_CSN   ;
wire        cap_FDA0_SDI   ;
wire        cap_DAC0_SCK   ;
wire        cap_DAC0_CSN   ;
wire        cap_DAC0_SDI   ;
wire        cap_OPA0_10X1  ;
wire        cap_OPA0_10X2  ;
wire        cap_OPA0_OPX1  ;
wire        cap_OPA0_OPX2  ;
Tc_PL_cap
#(
.TOP0_0     (TOP0_0     ),
.TOP0_1     (TOP0_1     ),
.TOP0_2     (TOP0_2     ),
.TOP0_3     (TOP0_3     ),
.TOP0_4     (TOP0_4     ),
.ADC0_0     (ADC0_0     ),
.ADC0_1     (ADC0_1     ),
.LDD0_0     (LDD0_0     ),
.CAP0_0     (CAP0_0     ),
.CAP0_1     (CAP0_1     ),
.AGP0_0     (AGP0_0     ),
.AGP0_1     (AGP0_1     ),
.AGP0_2     (AGP0_2     ),
.AGP0_3     (AGP0_3     ),
.AGP0_4     (AGP0_4     ),
.AGP0_5     (AGP0_5     ),
.AGP0_6     (AGP0_6     ),
.AGP0_7     (AGP0_7     ),
.AGP0_8     (AGP0_8     ),
.AGP0_9     (AGP0_9     ),
.AGP0_10    (AGP0_10    ),
.AGP0_11    (AGP0_11    ),
.AGP0_12    (AGP0_12    ),
.AGP0_13    (AGP0_13    ),
.AGP0_14    (AGP0_14    ),
.AGP0_15    (AGP0_15    ),
.AGP0_16    (AGP0_16    ),
.AGP0_17    (AGP0_17    ),
.AGP0_18    (AGP0_18    ),
.AGP0_19    (AGP0_19    ),
.AGP0_20    (AGP0_20    ),
.AGP0_21    (AGP0_21    ),
.AGP0_22    (AGP0_22    ),
.AGP0_23    (AGP0_23    ),
.AGP0_24    (AGP0_24    ),
.AGP0_25    (AGP0_25    ),
.AGP0_26    (AGP0_26    ),
.AGP0_27    (AGP0_27    ),
.AGP0_28    (AGP0_28    ),
.AGP0_29    (AGP0_29    ),
.AGP0_30    (AGP0_30    ),
.AGP0_31    (AGP0_31    ),
.AGP0_32    (AGP0_32    ),
.AGP0_33    (AGP0_33    ),
.AGP0_34    (AGP0_34    ),
.AGP0_35    (AGP0_35    )
)
Tc_PL_cap_ins0
(
.clk125           (clk125           ),
.rst              (rst              ),
.Gc_merge_data    (Gc_merge_data    ),
.Gc_mereg_datv    (Gc_mereg_datv    ),
.Gc_mereg_datr    (Gc_mereg_datr    ),
.Gc_cap_trig      (Gc_cap_trig      ),
.Gc_capr_rdy      (Gc_capr_rdy      ),
.Gc_cap_mode      (Gc_cap_mode      ),
.Gc_cap_wdis      (Gc_cap_wdis      ),
.Gc_cap_plus      (Gc_cap_plus      ),
.gp0_c0           (gp0_c0           ),
.gp0_c1           (gp0_c1           ),
.gp0_c2           (gp0_c2           ),
.gp0_c3           (gp0_c3           ),
.gp0_c4           (gp0_c4           ),
.gp0_c5           (gp0_c5           ),
.gp0_c6           (gp0_c6           ),
.gp0_c7           (gp0_c7           ),
.gp0_c8           (gp0_c8           ),
.gp0_c9           (gp0_c9           ),
.gp0_c10          (gp0_c10          ),
.gp0_c11          (gp0_c11          ),
.gp0_c12          (gp0_c12          ),
.gp0_c13          (gp0_c13          ),
.gp0_c14          (gp0_c14          ),
.gp0_c15          (gp0_c15          ),
.gp0_c16          (gp0_c16          ),
.gp0_c17          (gp0_c17          ),
.gp0_c18          (gp0_c18          ),
.gp0_c19          (gp0_c19          ),
.gp0_c20          (gp0_c20          ),
.gp0_c21          (gp0_c21          ),
.gp0_c22          (gp0_c22          ),
.gp0_c23          (gp0_c23          ),
.gp0_c24          (gp0_c24          ),
.gp0_c25          (gp0_c25          ),
.gp0_c26          (gp0_c26          ),
.gp0_c27          (gp0_c27          ),
.gp0_c28          (gp0_c28          ),
.gp0_c29          (gp0_c29          ),
.gp0_c30          (gp0_c30          ),
.gp0_c31          (gp0_c31          ),
.gp0_c32          (gp0_c32          ),
.gp0_c33          (gp0_c33          ),
.gp0_c34          (gp0_c34          ),
.gp0_c35          (gp0_c35          ),
.gp0_c0w          (gp0_c0w          ),
.acp0_tx_en       (acp0_tx_en       ),
.acp0_tx_rdy      (acp0_tx_rdy      ),
.acp0_tx_awaddr   (acp0_tx_awaddr   ),
.acp0_tx_awid     (acp0_tx_awid     ),
.acp0_tx_wdata    (acp0_tx_wdata    ),
.acp0_tx_wdreq    (acp0_tx_wdreq    ),
.FDA0_SCK         (cap_FDA0_SCK     ),
.FDA0_CSN         (cap_FDA0_CSN     ),
.FDA0_SDI         (cap_FDA0_SDI     ),
.DAC0_SDI         (cap_DAC0_SDI     ),
.DAC0_SCK         (cap_DAC0_SCK     ),
.DAC0_CSN         (cap_DAC0_CSN     ),
.OPA0_10X1        (cap_OPA0_10X1    ),
.OPA0_10X2        (cap_OPA0_10X2    ),
.OPA0_OPX1        (cap_OPA0_OPX1    ),
.OPA0_OPX2        (cap_OPA0_OPX2    )
    );

wire bus_FDA0_SCK;
wire bus_FDA0_CSN;
wire bus_FDA0_SDI;
wire bus_DAC0_SCK;
wire bus_DAC0_CSN;
wire bus_DAC0_SDI;
Tc_PL_bus
#(
.AGP0_21(AGP0_21	),
.AGP0_22(AGP0_22	),
.AGP0_23(AGP0_23	),
.AGP0_24(AGP0_24	),
.AGP0_25(AGP0_25	),
.AGP0_26(AGP0_26	),
.AGP0_27(AGP0_27	)
)
Tc_PL_bus_ins0
(
.clk         (clk125          ),
.rst         (rst             ),
.gp0_b0      (gp0_b0          ),
.gp0_b1      (gp0_b1          ),
.gp0_b2      (gp0_b2          ),
.gp0_b3      (gp0_b3          ),
.gp0_b4      (gp0_b4          ),
.gp0_b5      (gp0_b5          ),
.gp0_b6      (gp0_b6          ),
.gp0_b0w     (gp0_b0w         ),
.gp0_b2w     (gp0_b2w         ),
.gp0_b4r     (gp0_b4r         ),
.ADC0_CSN    (ADC0_CSN        ),
.ADC0_SCK    (ADC0_SCK        ),
.ADC0_SDI    (ADC0_SDI        ),
.ADC0_SDO    (ADC0_SDO        ),
.FDA0_SCK    (bus_FDA0_SCK    ),
.FDA0_CSN    (bus_FDA0_CSN    ),
.FDA0_SDI    (bus_FDA0_SDI    ),
.FDA0_SDO    (FDA0_SDO        ),
.DAC0_SDI    (bus_DAC0_SDI    ),
.DAC0_SCK    (bus_DAC0_SCK    ),
.DAC0_CSN    (bus_DAC0_CSN    ),
.DAC1_SDI    (DAC1_SDI        ),
.DAC1_SCK    (DAC1_SCK        ),
.DAC1_CSN    (DAC1_CSN        ),
.LPL0_CSN    (LPL0_CSN        ),
.LPL0_SDO    (LPL0_SDO        ),
.LPL0_SCK    (LPL0_SCK        ),
.LPL0_SDI    (LPL0_SDI        )
    );

wire                   chips_OPA0_10X1 ;
wire                   chips_OPA0_10X2 ;
wire                   chips_OPA0_OPX1 ;
wire                   chips_OPA0_OPX2 ;
Tc_PL_chips
#(
.TOP0_0    (TOP0_0    ),
.TOP0_1    (TOP0_1    ),
.TOP0_2    (TOP0_2    ),
.TOP0_3    (TOP0_3    ),
.TOP0_4    (TOP0_4    ),
.ADC0_0    (ADC0_0    ),
.ADC0_1    (ADC0_1    ),
.LDD0_0    (LDD0_0    ),
.CAP0_0    (CAP0_0    ),
.CAP0_1    (CAP0_1    ),
.AGP0_0    (AGP0_0    ),
.AGP0_1    (AGP0_1    ),
.AGP0_2    (AGP0_2    ),
.AGP0_3    (AGP0_3    ),
.AGP0_4    (AGP0_4    ),
.AGP0_5    (AGP0_5    ),
.AGP0_6    (AGP0_6    ),
.AGP0_7    (AGP0_7    ),
.AGP0_8    (AGP0_8    ),
.AGP0_9    (AGP0_9    ),
.AGP0_10   (AGP0_10   ),
.AGP0_11   (AGP0_11   ),
.AGP0_12   (AGP0_12   ),
.AGP0_13   (AGP0_13   ),
.AGP0_14   (AGP0_14   ),
.AGP0_15   (AGP0_15   ),
.AGP0_16   (AGP0_16   ),
.AGP0_17   (AGP0_17   ),
.AGP0_18   (AGP0_18   ),
.AGP0_19   (AGP0_19   ),
.AGP0_20   (AGP0_20   ),
.AGP0_21   (AGP0_21   ),
.AGP0_22   (AGP0_22   ),
.AGP0_23   (AGP0_23   ),
.AGP0_24   (AGP0_24   ),
.AGP0_25   (AGP0_25   ),
.AGP0_26   (AGP0_26   ),
.AGP0_27   (AGP0_27   ),
.AGP0_28   (AGP0_28   ),
.AGP0_29   (AGP0_29   ),
.AGP0_30   (AGP0_30   ),
.AGP0_31   (AGP0_31   ),
.AGP0_32   (AGP0_32   ),
.AGP0_33   (AGP0_33   ),
.AGP0_34   (AGP0_34   ),
.AGP0_35   (AGP0_35   )
)
Tc_PL_chips_ins0
(
.clk125        (clk125        ),
.rst           (rst           ),
.Gc_adc_of     (Gc_adc_of     ),
.Gc_adc_data   (Gc_adc_data   ),
.Gc_com_wdis   (Gc_com_wdis   ),
.Gc_com_plus   (Gc_com_plus   ),
.Gc_com_open   (Gc_com_open   ),
.Gc_com_close  (Gc_com_close  ),
.Gc_wdis       (Gc_wdis       ),
.gp0_d0        (gp0_d0        ),
.gp0_d1        (gp0_d1        ),
.gp0_d2        (gp0_d2        ),
.gp0_d3        (gp0_d3        ),
.gp0_d4        (gp0_d4        ),
.gp0_d5        (gp0_d5        ),
.gp0_r0        (gp0_r0        ),
.gp0_r1        (gp0_r1        ),
.gp0_r2        (gp0_r2        ),
.gp0_r3        (gp0_r3        ),
.gp0_r4        (gp0_r4        ),
.gp0_r5        (gp0_r5        ),
.gp0_r6        (gp0_r6        ),
.gp0_r7        (gp0_r7        ),
.gp0_r7w       (gp0_r7w       ),
.LDD0_OUTEA    (LDD0_OUTEA    ),
.LDD0_DISEA    (LDD0_DISEA    ),
.LDD0_OSCEA    (LDD0_OSCEA    ),
.LDD0_OLD2N    (LDD0_OLD2N    ),
.LDD0_RDISN    (LDD0_RDISN    ),
.OPA0_10X1     (chips_OPA0_10X1     ),
.OPA0_10X2     (chips_OPA0_10X2     ),
.OPA0_OPX1     (chips_OPA0_OPX1     ),
.OPA0_OPX2     (chips_OPA0_OPX2     ),
.APD0_EN       (APD0_EN       ),
.LPL0_LOCK     (LPL0_LOCK     ),
.LPL0_ERR      (LPL0_ERR      ),
.LPL0_SYNC     (LPL0_SYNC     ),
.TEC0_GOOD     (TEC0_GOOD     ),
.TEC1_GOOD     (TEC1_GOOD     ),
.LED0_L        (LED0_L        ),
.OPM0_IO       (OPM0_IO       )
    );

assign FDA0_SCK  = Gc_cap_mode ? cap_FDA0_SCK : bus_FDA0_SCK   ;
assign FDA0_CSN  = Gc_cap_mode ? cap_FDA0_CSN : bus_FDA0_CSN   ;
assign FDA0_SDI  = Gc_cap_mode ? cap_FDA0_SDI : bus_FDA0_SDI   ;
assign DAC0_SCK  = Gc_cap_mode ? cap_DAC0_SCK : bus_DAC0_SCK   ;
assign DAC0_CSN  = Gc_cap_mode ? cap_DAC0_CSN : bus_DAC0_CSN   ;
assign DAC0_SDI  = Gc_cap_mode ? cap_DAC0_SDI : bus_DAC0_SDI   ;
assign OPA0_10X1 = Gc_cap_mode ? cap_OPA0_10X1: chips_OPA0_10X1;
assign OPA0_10X2 = Gc_cap_mode ? cap_OPA0_10X2: chips_OPA0_10X2;
assign OPA0_OPX1 = Gc_cap_mode ? cap_OPA0_OPX1: chips_OPA0_OPX1;
assign OPA0_OPX2 = Gc_cap_mode ? cap_OPA0_OPX2: chips_OPA0_OPX2;

endmodule
