`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2020/02/09 12:20:59
// Design Name:
// Module Name: Tc_PS_Zynq
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module Tc_PS_Zynq(
inout      [14:0]     DDR_addr                 ,
inout      [2:0]      DDR_ba                   ,
inout                 DDR_cas_n                ,
inout                 DDR_ck_n                 ,
inout                 DDR_ck_p                 ,
inout                 DDR_cke                  ,
inout                 DDR_cs_n                 ,
inout      [3:0]      DDR_dm                   ,
inout      [31:0]     DDR_dq                   ,
inout      [3:0]      DDR_dqs_n                ,
inout      [3:0]      DDR_dqs_p                ,
inout                 DDR_odt                  ,
inout                 DDR_ras_n                ,
inout                 DDR_reset_n              ,
inout                 DDR_we_n                 ,
output                FCLK_CLK0_0              ,
output                FCLK_RESET0_N_0          ,
inout                 FIXED_IO_ddr_vrn         ,
inout                 FIXED_IO_ddr_vrp         ,
inout      [53:0]     FIXED_IO_mio             ,
inout                 FIXED_IO_ps_clk          ,
inout                 FIXED_IO_ps_porb         ,
inout                 FIXED_IO_ps_srstb        ,
input      [63:0]     GPIO_I_0                 ,
output     [63:0]     GPIO_O_0                 ,
output     [63:0]     GPIO_T_0                 ,
input      [15:0]     IRQ_F2P_0                ,
output     [31:0]     M_AXI_GP0_0_araddr       ,
output     [1:0]      M_AXI_GP0_0_arburst      ,
output     [3:0]      M_AXI_GP0_0_arcache      ,
output     [11:0]     M_AXI_GP0_0_arid         ,
output     [3:0]      M_AXI_GP0_0_arlen        ,
output     [1:0]      M_AXI_GP0_0_arlock       ,
output     [2:0]      M_AXI_GP0_0_arprot       ,
output     [3:0]      M_AXI_GP0_0_arqos        ,
input                 M_AXI_GP0_0_arready      ,
output     [2:0]      M_AXI_GP0_0_arsize       ,
output                M_AXI_GP0_0_arvalid      ,
output     [31:0]     M_AXI_GP0_0_awaddr       ,
output     [1:0]      M_AXI_GP0_0_awburst      ,
output     [3:0]      M_AXI_GP0_0_awcache      ,
output     [11:0]     M_AXI_GP0_0_awid         ,
output     [3:0]      M_AXI_GP0_0_awlen        ,
output     [1:0]      M_AXI_GP0_0_awlock       ,
output     [2:0]      M_AXI_GP0_0_awprot       ,
output     [3:0]      M_AXI_GP0_0_awqos        ,
input                 M_AXI_GP0_0_awready      ,
output     [2:0]      M_AXI_GP0_0_awsize       ,
output                M_AXI_GP0_0_awvalid      ,
input      [11:0]     M_AXI_GP0_0_bid          ,
output                M_AXI_GP0_0_bready       ,
input      [1:0]      M_AXI_GP0_0_bresp        ,
input                 M_AXI_GP0_0_bvalid       ,
input      [31:0]     M_AXI_GP0_0_rdata        ,
input      [11:0]     M_AXI_GP0_0_rid          ,
input                 M_AXI_GP0_0_rlast        ,
output                M_AXI_GP0_0_rready       ,
input      [1:0]      M_AXI_GP0_0_rresp        ,
input                 M_AXI_GP0_0_rvalid       ,
output     [31:0]     M_AXI_GP0_0_wdata        ,
output     [11:0]     M_AXI_GP0_0_wid          ,
output                M_AXI_GP0_0_wlast        ,
input                 M_AXI_GP0_0_wready       ,
output     [3:0]      M_AXI_GP0_0_wstrb        ,
output                M_AXI_GP0_0_wvalid       ,
input                 M_AXI_GP0_ACLK_0         ,
input                 SPI0_MISO_I_0            ,
output                SPI0_MOSI_O_0            ,
output                SPI0_SCLK_O_0            ,
output                SPI0_SS1_O_0             ,
output                SPI0_SS2_O_0             ,
output                SPI0_SS_O_0              ,
input      [31:0]     S_AXI_ACP_0_araddr       ,
input      [1:0]      S_AXI_ACP_0_arburst      ,
input      [3:0]      S_AXI_ACP_0_arcache      ,
input      [2:0]      S_AXI_ACP_0_arid         ,
input      [3:0]      S_AXI_ACP_0_arlen        ,
input      [1:0]      S_AXI_ACP_0_arlock       ,
input      [2:0]      S_AXI_ACP_0_arprot       ,
input      [3:0]      S_AXI_ACP_0_arqos        ,
output                S_AXI_ACP_0_arready      ,
input      [2:0]      S_AXI_ACP_0_arsize       ,
input      [4:0]      S_AXI_ACP_0_aruser       ,
input                 S_AXI_ACP_0_arvalid      ,
input      [31:0]     S_AXI_ACP_0_awaddr       ,
input      [1:0]      S_AXI_ACP_0_awburst      ,
input      [3:0]      S_AXI_ACP_0_awcache      ,
input      [2:0]      S_AXI_ACP_0_awid         ,
input      [3:0]      S_AXI_ACP_0_awlen        ,
input      [1:0]      S_AXI_ACP_0_awlock       ,
input      [2:0]      S_AXI_ACP_0_awprot       ,
input      [3:0]      S_AXI_ACP_0_awqos        ,
output                S_AXI_ACP_0_awready      ,
input      [2:0]      S_AXI_ACP_0_awsize       ,
input      [4:0]      S_AXI_ACP_0_awuser       ,
input                 S_AXI_ACP_0_awvalid      ,
output     [2:0]      S_AXI_ACP_0_bid          ,
input                 S_AXI_ACP_0_bready       ,
output     [1:0]      S_AXI_ACP_0_bresp        ,
output                S_AXI_ACP_0_bvalid       ,
output     [63:0]     S_AXI_ACP_0_rdata        ,
output     [2:0]      S_AXI_ACP_0_rid          ,
output                S_AXI_ACP_0_rlast        ,
input                 S_AXI_ACP_0_rready       ,
output     [1:0]      S_AXI_ACP_0_rresp        ,
output                S_AXI_ACP_0_rvalid       ,
input      [63:0]     S_AXI_ACP_0_wdata        ,
input      [2:0]      S_AXI_ACP_0_wid          ,
input                 S_AXI_ACP_0_wlast        ,
output                S_AXI_ACP_0_wready       ,
input      [7:0]      S_AXI_ACP_0_wstrb        ,
input                 S_AXI_ACP_0_wvalid       ,
input                 S_AXI_ACP_ACLK_0         ,
input                 UART_0_0_rxd             ,
output                UART_0_0_txd
    );

IRLv2_wrapper
IRLv2_wrapper_ins0
(
.DDR_addr            (DDR_addr                   ),
.DDR_ba              (DDR_ba                     ),
.DDR_cas_n           (DDR_cas_n                  ),
.DDR_ck_n            (DDR_ck_n                   ),
.DDR_ck_p            (DDR_ck_p                   ),
.DDR_cke             (DDR_cke                    ),
.DDR_cs_n            (DDR_cs_n                   ),
.DDR_dm              (DDR_dm                     ),
.DDR_dq              (DDR_dq                     ),
.DDR_dqs_n           (DDR_dqs_n                  ),
.DDR_dqs_p           (DDR_dqs_p                  ),
.DDR_odt             (DDR_odt                    ),
.DDR_ras_n           (DDR_ras_n                  ),
.DDR_reset_n         (DDR_reset_n                ),
.DDR_we_n            (DDR_we_n                   ),
.FCLK_CLK0_0         (FCLK_CLK0_0                ),
.FCLK_RESET0_N_0     (FCLK_RESET0_N_0            ),
.FIXED_IO_ddr_vrn    (FIXED_IO_ddr_vrn           ),
.FIXED_IO_ddr_vrp    (FIXED_IO_ddr_vrp           ),
.FIXED_IO_mio        (FIXED_IO_mio               ),
.FIXED_IO_ps_clk     (FIXED_IO_ps_clk            ),
.FIXED_IO_ps_porb    (FIXED_IO_ps_porb           ),
.FIXED_IO_ps_srstb   (FIXED_IO_ps_srstb          ),
.GPIO_I_0            (GPIO_I_0                   ),
.GPIO_O_0            (GPIO_O_0                   ),
.GPIO_T_0            (GPIO_T_0                   ),
.IRQ_F2P_0           (IRQ_F2P_0                  ),
.M_AXI_GP0_0_araddr  (M_AXI_GP0_0_araddr         ),
.M_AXI_GP0_0_arburst (M_AXI_GP0_0_arburst        ),
.M_AXI_GP0_0_arcache (M_AXI_GP0_0_arcache        ),
.M_AXI_GP0_0_arid    (M_AXI_GP0_0_arid           ),
.M_AXI_GP0_0_arlen   (M_AXI_GP0_0_arlen          ),
.M_AXI_GP0_0_arlock  (M_AXI_GP0_0_arlock         ),
.M_AXI_GP0_0_arprot  (M_AXI_GP0_0_arprot         ),
.M_AXI_GP0_0_arqos   (M_AXI_GP0_0_arqos          ),
.M_AXI_GP0_0_arready (M_AXI_GP0_0_arready        ),
.M_AXI_GP0_0_arsize  (M_AXI_GP0_0_arsize         ),
.M_AXI_GP0_0_arvalid (M_AXI_GP0_0_arvalid        ),
.M_AXI_GP0_0_awaddr  (M_AXI_GP0_0_awaddr         ),
.M_AXI_GP0_0_awburst (M_AXI_GP0_0_awburst        ),
.M_AXI_GP0_0_awcache (M_AXI_GP0_0_awcache        ),
.M_AXI_GP0_0_awid    (M_AXI_GP0_0_awid           ),
.M_AXI_GP0_0_awlen   (M_AXI_GP0_0_awlen          ),
.M_AXI_GP0_0_awlock  (M_AXI_GP0_0_awlock         ),
.M_AXI_GP0_0_awprot  (M_AXI_GP0_0_awprot         ),
.M_AXI_GP0_0_awqos   (M_AXI_GP0_0_awqos          ),
.M_AXI_GP0_0_awready (M_AXI_GP0_0_awready        ),
.M_AXI_GP0_0_awsize  (M_AXI_GP0_0_awsize         ),
.M_AXI_GP0_0_awvalid (M_AXI_GP0_0_awvalid        ),
.M_AXI_GP0_0_bid     (M_AXI_GP0_0_bid            ),
.M_AXI_GP0_0_bready  (M_AXI_GP0_0_bready         ),
.M_AXI_GP0_0_bresp   (M_AXI_GP0_0_bresp          ),
.M_AXI_GP0_0_bvalid  (M_AXI_GP0_0_bvalid         ),
.M_AXI_GP0_0_rdata   (M_AXI_GP0_0_rdata          ),
.M_AXI_GP0_0_rid     (M_AXI_GP0_0_rid            ),
.M_AXI_GP0_0_rlast   (M_AXI_GP0_0_rlast          ),
.M_AXI_GP0_0_rready  (M_AXI_GP0_0_rready         ),
.M_AXI_GP0_0_rresp   (M_AXI_GP0_0_rresp          ),
.M_AXI_GP0_0_rvalid  (M_AXI_GP0_0_rvalid         ),
.M_AXI_GP0_0_wdata   (M_AXI_GP0_0_wdata          ),
.M_AXI_GP0_0_wid     (M_AXI_GP0_0_wid            ),
.M_AXI_GP0_0_wlast   (M_AXI_GP0_0_wlast          ),
.M_AXI_GP0_0_wready  (M_AXI_GP0_0_wready         ),
.M_AXI_GP0_0_wstrb   (M_AXI_GP0_0_wstrb          ),
.M_AXI_GP0_0_wvalid  (M_AXI_GP0_0_wvalid         ),
.M_AXI_GP0_ACLK_0    (M_AXI_GP0_ACLK_0           ),
.SPI0_MISO_I_0       (SPI0_MISO_I_0              ),
.SPI0_MOSI_O_0       (SPI0_MOSI_O_0              ),
.SPI0_SCLK_O_0       (SPI0_SCLK_O_0              ),
.SPI0_SS1_O_0        (SPI0_SS1_O_0               ),
.SPI0_SS2_O_0        (SPI0_SS2_O_0               ),
.SPI0_SS_O_0         (SPI0_SS_O_0                ),
.S_AXI_ACP_0_araddr  (S_AXI_ACP_0_araddr         ),
.S_AXI_ACP_0_arburst (S_AXI_ACP_0_arburst        ),
.S_AXI_ACP_0_arcache (S_AXI_ACP_0_arcache        ),
.S_AXI_ACP_0_arid    (S_AXI_ACP_0_arid           ),
.S_AXI_ACP_0_arlen   (S_AXI_ACP_0_arlen          ),
.S_AXI_ACP_0_arlock  (S_AXI_ACP_0_arlock         ),
.S_AXI_ACP_0_arprot  (S_AXI_ACP_0_arprot         ),
.S_AXI_ACP_0_arqos   (S_AXI_ACP_0_arqos          ),
.S_AXI_ACP_0_arready (S_AXI_ACP_0_arready        ),
.S_AXI_ACP_0_arsize  (S_AXI_ACP_0_arsize         ),
.S_AXI_ACP_0_aruser  (S_AXI_ACP_0_aruser         ),
.S_AXI_ACP_0_arvalid (S_AXI_ACP_0_arvalid        ),
.S_AXI_ACP_0_awaddr  (S_AXI_ACP_0_awaddr         ),
.S_AXI_ACP_0_awburst (S_AXI_ACP_0_awburst        ),
.S_AXI_ACP_0_awcache (S_AXI_ACP_0_awcache        ),
.S_AXI_ACP_0_awid    (S_AXI_ACP_0_awid           ),
.S_AXI_ACP_0_awlen   (S_AXI_ACP_0_awlen          ),
.S_AXI_ACP_0_awlock  (S_AXI_ACP_0_awlock         ),
.S_AXI_ACP_0_awprot  (S_AXI_ACP_0_awprot         ),
.S_AXI_ACP_0_awqos   (S_AXI_ACP_0_awqos          ),
.S_AXI_ACP_0_awready (S_AXI_ACP_0_awready        ),
.S_AXI_ACP_0_awsize  (S_AXI_ACP_0_awsize         ),
.S_AXI_ACP_0_awuser  (S_AXI_ACP_0_awuser         ),
.S_AXI_ACP_0_awvalid (S_AXI_ACP_0_awvalid        ),
.S_AXI_ACP_0_bid     (S_AXI_ACP_0_bid            ),
.S_AXI_ACP_0_bready  (S_AXI_ACP_0_bready         ),
.S_AXI_ACP_0_bresp   (S_AXI_ACP_0_bresp          ),
.S_AXI_ACP_0_bvalid  (S_AXI_ACP_0_bvalid         ),
.S_AXI_ACP_0_rdata   (S_AXI_ACP_0_rdata          ),
.S_AXI_ACP_0_rid     (S_AXI_ACP_0_rid            ),
.S_AXI_ACP_0_rlast   (S_AXI_ACP_0_rlast          ),
.S_AXI_ACP_0_rready  (S_AXI_ACP_0_rready         ),
.S_AXI_ACP_0_rresp   (S_AXI_ACP_0_rresp          ),
.S_AXI_ACP_0_rvalid  (S_AXI_ACP_0_rvalid         ),
.S_AXI_ACP_0_wdata   (S_AXI_ACP_0_wdata          ),
.S_AXI_ACP_0_wid     (S_AXI_ACP_0_wid            ),
.S_AXI_ACP_0_wlast   (S_AXI_ACP_0_wlast          ),
.S_AXI_ACP_0_wready  (S_AXI_ACP_0_wready         ),
.S_AXI_ACP_0_wstrb   (S_AXI_ACP_0_wstrb          ),
.S_AXI_ACP_0_wvalid  (S_AXI_ACP_0_wvalid         ),
.S_AXI_ACP_ACLK_0    (S_AXI_ACP_ACLK_0           ),
.UART_0_0_rxd        (UART_0_0_rxd               ),
.UART_0_0_txd        (UART_0_0_txd               )
);

endmodule
